package shared_pkg;
bit test_finished;
int error_count;
int correct_count;
event etrigger;
endpackage

